
module Internal_OSC (
	oscena,
	clkout);	

	input		oscena;
	output		clkout;
endmodule
