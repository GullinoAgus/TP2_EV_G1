// megafunction wizard: %ALTDDIO_IN%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTDDIO_IN 

// ============================================================
// File Name: pin_io.v
// Megafunction Name(s):
// 			ALTDDIO_IN
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 23.1std.0 Build 991 11/28/2023 SC Lite Edition
// ************************************************************

//Copyright (C) 2023  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and any partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details, at
//https://fpgasoftware.intel.com/eula.

module pin_io (
	datain,
	inclock,
	dataout_h,
	dataout_l);

	input	[31:0]  datain;
	input	  inclock;
	output	[31:0]  dataout_h;
	output	[31:0]  dataout_l;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: CONSTANT: INVERT_INPUT_CLOCKS STRING "OFF"
// Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altddio_in"
// Retrieval info: CONSTANT: POWER_UP_HIGH STRING "OFF"
// Retrieval info: CONSTANT: WIDTH NUMERIC "32"
// Retrieval info: USED_PORT: datain 0 0 32 0 INPUT NODEFVAL "datain[31..0]"
// Retrieval info: CONNECT: @datain 0 0 32 0 datain 0 0 32 0
// Retrieval info: USED_PORT: dataout_h 0 0 32 0 OUTPUT NODEFVAL "dataout_h[31..0]"
// Retrieval info: CONNECT: dataout_h 0 0 32 0 @dataout_h 0 0 32 0
// Retrieval info: USED_PORT: dataout_l 0 0 32 0 OUTPUT NODEFVAL "dataout_l[31..0]"
// Retrieval info: CONNECT: dataout_l 0 0 32 0 @dataout_l 0 0 32 0
// Retrieval info: USED_PORT: inclock 0 0 0 0 INPUT_CLK_EXT NODEFVAL "inclock"
// Retrieval info: CONNECT: @inclock 0 0 0 0 inclock 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL pin_io.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL pin_io.qip TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL pin_io.bsf TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL pin_io_inst.v FALSE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL pin_io_bb.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL pin_io.inc FALSE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL pin_io.cmp FALSE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL pin_io.ppf TRUE FALSE
// Retrieval info: LIB_FILE: altera_mf
