module decode(

);


endmodule